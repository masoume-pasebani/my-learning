
module ALU( out_put , A , B ,sel);
  output out_put;
  input A;
  input B;
  input sel;
endmodule
