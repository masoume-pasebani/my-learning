
module ALU( out_put , A , B ,sel,co);
  output out_put;
  input [7:0] A;
  input [7:0] B;
  input [1:0] sel;
endmodule
