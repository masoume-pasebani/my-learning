module operation_0();
endmodule
